`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.08.2020 20:16:50
// Design Name: 
// Module Name: mips_test
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mips_test( );
reg clk1,clk2;
integer k;

Mips mips (clk1,clk2);

initial
    begin
        clk1=0;clk2=0;
        repeat(50)
        begin
            #5 clk1=1; 
            #5 clk1=0;
            #5 clk2=1;
            #5 clk2=1;
        end
    end
    
    initial
        begin
            for(k=0;k<31;k=k+1)
            mips.Reg[k]=k;
            
            mips.Mem[0] =32'h280a00c8; //ADDI R10,R0,200
            mips.Mem[1] = 32'h28020001;//ADDI R2,R0,1
            mips.Mem[2]=32'h0e94a000;//OR R20,R20,R20 --- DUMMT
            mips.Mem[3] = 32'h21430000;//LW R3,0(R10)
            mips.Mem[4] = 32'h0e94a000;//OR R20,R20,20  --DUMY
            mips.Mem[5] = 32'h14431000;//LOOP MUL R2,R2,R3
            mips.Mem[6] = 32'h2c630001;//SUBI R3,R3,1
            mips.Mem[7] = 32'h0e94a000;//OR R20,R20,R20
            mips.Mem[8] = 32'h3460fffc;//BNEQZ R3,LOOP
            mips.Mem[9] = 32'h2542fffe;//SW R2.-2(R10)
            mips.Mem[10] = 32'hfc000000;//HLT
            
            mips.HALTED =0;
            mips.PC=0;
            mips.TAKEN_BRANCH =0;
            
            #300
            for(k=0;k<6;k=k+1)
            $dispay("R%1d -%2d", k, mips.Reg[k]);
            //#300 finish;
        end
endmodule
